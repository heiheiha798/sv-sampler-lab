module component_0(
    input wire [28:0] var_0,
    input wire [26:0] var_1,
    input wire [12:0] var_2,
    input wire [23:0] var_3,
    input wire [3:0] var_4,
    input wire [9:0] var_6,
    input wire [16:0] var_7,
    input wire [11:0] var_8,
    input wire [31:0] var_9,
    input wire [20:0] var_11,
    input wire [13:0] var_12,
    input wire [31:0] var_13,
    input wire [7:0] var_14,
    input wire [17:0] var_15,
    input wire [7:0] var_16,
    input wire [17:0] var_18,
    input wire [8:0] var_20,
    input wire [17:0] var_21,
    input wire [10:0] var_22,
    input wire [3:0] var_23,
    input wire [6:0] var_24,
    input wire [29:0] var_25,
    input wire [26:0] var_26,
    input wire [26:0] var_28,
    input wire [6:0] var_29,
    output wire result
);

    wire cnstr_1_w;
    wire cnstr_2_w;
    wire cnstr_0_w;
    wire cnstr_3_w;
    wire cnstr_4_w;
    wire cnstr_5_w;
    wire cnstr_7_w;
    wire cnstr_8_w;
    wire cnstr_9_w;
    wire cnstr_10_w;
    wire cnstr_11_w;
    wire cnstr_12_w;
    wire cnstr_15_w;
    wire cnstr_17_w;
    wire cnstr_18_w;
    wire cnstr_19_w;
    wire cnstr_20_w;
    wire cnstr_21_w;
    wire cnstr_22_w;
    wire cnstr_23_w;
    wire cnstr_24_w;
    wire cnstr_25_w;
    wire cnstr_26_w;
    wire cnstr_28_w;
    wire cnstr_29_w;
    wire cnstr_6_w;
    wire cnstr_13_w;
    wire cnstr_14_w;
    wire cnstr_16_w;
    wire cnstr_27_w;

    assign cnstr_1_w = |(~((var_11 + 32'h853b9)));
    assign cnstr_2_w = |((var_2 | 13'h19de));
    assign cnstr_0_w = |((var_14 * var_29));
    assign cnstr_3_w = |(( (!(var_24)) || (var_29) ));
    assign cnstr_4_w = |((var_0 || var_3));
    assign cnstr_5_w = |(((var_7 & var_4) != var_18));
    assign cnstr_7_w = |((var_28 - var_14));
    assign cnstr_8_w = |(( (!(var_21)) || (var_4) ));
    assign cnstr_9_w = |((~(var_25) | var_1));
    assign cnstr_10_w = |(((var_16 / 8'h4) && var_6));
    assign cnstr_11_w = |(((var_16 * var_14) != var_21));
    assign cnstr_12_w = |(!((var_0 + var_26)));
    assign cnstr_15_w = |(((var_22 + 32'h41e) - 32'h276a248e));
    assign cnstr_17_w = |((var_26 != var_15));
    assign cnstr_18_w = |(~((var_21 && var_25)));
    assign cnstr_19_w = |(!(~((var_24 * 8'h5))));
    assign cnstr_20_w = |((~(var_21) << 18'h1));
    assign cnstr_21_w = |((var_26 << 27'h6));
    assign cnstr_22_w = |((var_20 | var_24));
    assign cnstr_23_w = |((!(var_8) || var_29));
    assign cnstr_24_w = |((var_21 << 18'h0));
    assign cnstr_25_w = |((var_25 || var_6));
    assign cnstr_26_w = |(!((var_4 + var_26)));
    assign cnstr_28_w = |(((var_1 | var_22) | var_16));
    assign cnstr_29_w = |((var_14 != 32'hb8));
    assign cnstr_6_w = |((var_12 | 14'h2cd9));
    assign cnstr_13_w = |(!((var_13 + 32'h75f0b4e2)));
    assign cnstr_14_w = |((~(var_23) / 4'h7));
    assign cnstr_16_w = |(( (!(var_9)) || (32'h6fbe9481) ));
    assign cnstr_27_w = |((var_9 ^ 32'h6839a06f));

    assign result = cnstr_1_w & cnstr_2_w & cnstr_6_w & cnstr_13_w & cnstr_14_w & cnstr_16_w & cnstr_27_w & cnstr_0_w & cnstr_3_w & cnstr_4_w & cnstr_5_w & cnstr_7_w & cnstr_8_w & cnstr_9_w & cnstr_10_w & cnstr_11_w & cnstr_12_w & cnstr_15_w & cnstr_17_w & cnstr_18_w & cnstr_19_w & cnstr_20_w & cnstr_21_w & cnstr_22_w & cnstr_23_w & cnstr_24_w & cnstr_25_w & cnstr_26_w & cnstr_28_w & cnstr_29_w;
endmodule
